module addOne
(
    input wire [4:0] I,
    output wire [4:0] O
);
assign O = I + 1;
endmodule